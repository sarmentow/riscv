module insmem(address, ins_out);
	input [31:0] address;
	output [31:0] ins_out;

	// 100 32 bit instruction capacity = 400 1 byte pieces of
	// instruction
	reg [7:0] ins [399:0];

	integer i;
	initial begin
		for (i = 0; i < 400; i = i + 1) begin
			ins[i] = 32'b0;
		end
		// addi x1, x0, 2
		ins[0] <= 8'b10010011;
		ins[1] <= 8'b00000000;
		ins[2] <= 8'b00100000;
		ins[3] <= 8'b00000000;

		// sw x1, 0(x0)
		ins[4] <= 8'b00100011;
		ins[5] <= 8'b00100000;
		ins[6] <= 8'b00010000;
		ins[7] <= 8'b00000000;

		// addi x1, x0, 3
		ins[8] <= 8'b10010011;
		ins[9] <= 8'b00000000;
		ins[10] <= 8'b00110000;
		ins[11] <= 8'b00000000;

		// sw x1, 4(x0)
		ins[12] <= 8'b00100011;
		ins[13] <= 8'b00100010;
		ins[14] <= 8'b00010000;
		ins[15] <= 8'b00000000;

		// addi x1, x0, 4
		ins[16] <= 8'b10010011;
		ins[17] <= 8'b00000000;
		ins[18] <= 8'b01000000;
		ins[19] <= 8'b00000000;

		// sw x1, 8(x0)
		ins[20] <= 8'b00100011;
		ins[21] <= 8'b00100100;
		ins[22] <= 8'b00010000;
		ins[23] <= 8'b00000000;

		// addi x1, x0, 8
		ins[24] <= 8'b10010011;
		ins[25] <= 8'b00000000;
		ins[26] <= 8'b10000000;
		ins[27] <= 8'b00000000;

		// sw x1, 12(x0)
		ins[28] <= 8'b00100011;
		ins[29] <= 8'b00100110;
		ins[30] <= 8'b00010000;
		ins[31] <= 8'b00000000;

		// addi x1, x0, 21
		ins[32] <= 8'b10010011;
		ins[33] <= 8'b00000000;
		ins[34] <= 8'b01010000;
		ins[35] <= 8'b00000001;

		// sw x1, 16(x0)
		ins[36] <= 8'b00100011;
		ins[37] <= 8'b00101000;
		ins[38] <= 8'b00010000;
		ins[39] <= 8'b00000000;

		// addi x1, x0, 2 
		ins[40] <= 8'b10010011;
		ins[41] <= 8'b00000000;
		ins[42] <= 8'b00100000;
		ins[43] <= 8'b00000000;

		// sw x1, 20(x0)
		ins[44] <= 8'b00100011;
		ins[45] <= 8'b00101010;
		ins[46] <= 8'b00010000;
		ins[47] <= 8'b00000000;

		// addi x1, x0, 30
		ins[48] <= 8'b10010011;
		ins[49] <= 8'b00000000;
		ins[50] <= 8'b11100000;
		ins[51] <= 8'b00000001;

		// sw x1, 24(x0)
		ins[52] <= 8'b00100011;
		ins[53] <= 8'b00101100;
		ins[54] <= 8'b00010000;
		ins[55] <= 8'b00000000;

		// addi x1, x0, 100
		ins[56] <= 8'b10010011;
		ins[57] <= 8'b00000000;
		ins[58] <= 8'b01000000;
		ins[59] <= 8'b00000110;

		// sw x1, 28(x0)
		ins[60] <= 8'b00100011;
		ins[61] <= 8'b00101110;
		ins[62] <= 8'b00010000;
		ins[63] <= 8'b00000000;

		// addi x1, x0, 31
		ins[64] <= 8'b10010011;
		ins[65] <= 8'b00000000;
		ins[66] <= 8'b11110000;
		ins[67] <= 8'b00000001;

		// sw x1, 32(x0)
		ins[68] <= 8'b00100011;
		ins[69] <= 8'b00100000;
		ins[70] <= 8'b00010000;
		ins[71] <= 8'b00000010;

		// addi x1, x0, 36
		ins[72] <= 8'b10010011;
		ins[73] <= 8'b00000000;
		ins[74] <= 8'b01000000;
		ins[75] <= 8'b00000010;

		// addi x2, x0, 0
		ins[76] <= 8'b00010011;
		ins[77] <= 8'b00000001;
		ins[78] <= 8'b00000000;
		ins[79] <= 8'b00000000;

		// lw x3, 0(x2)
		ins[80] <= 8'b10000011;
		ins[81] <= 8'b00100001;
		ins[82] <= 8'b00000001;
		ins[83] <= 8'b00000000;

		// bge x2, x1, 28 
		ins[84] <= 8'b01100011;
		ins[85] <= 8'b01011110;
		ins[86] <= 8'b00010001;
		ins[87] <= 8'b00000000;

		// lw x4, 0(x2)
		ins[88] <= 8'b00000011;
		ins[89] <= 8'b00100010;
		ins[90] <= 8'b00000001;
		ins[91] <= 8'b00000000;

		// addi x0, x0, 0
		ins[92] <= 8'b00010011;
		ins[93] <= 8'b00000000;
		ins[94] <= 8'b00000000;
		ins[95] <= 8'b00000000;

		// bge x3, x4, 8
		ins[96] <= 8'b01100011;
		ins[97] <= 8'b11010100;
		ins[98] <= 8'b01000001;
		ins[99] <= 8'b00000000;

		// add x3, x4, x0
		ins[100] <= 8'b10110011;
		ins[101] <= 8'b00000001;
		ins[102] <= 8'b00000010;
		ins[103] <= 8'b00000000;

		// addi x2, x2, 4
		ins[104] <= 8'b00010011;
		ins[105] <= 8'b00000001;
		ins[106] <= 8'b01000001;
		ins[107] <= 8'b00000000;

		// jal x0, -24
		ins[108] <= 8'b01101111;
		ins[109] <= 8'b11110000;
		ins[110] <= 8'b10011111;
		ins[111] <= 8'b11111110;

		// addi x0, x0, 0
		ins[112] <= 8'b00010011;
		ins[113] <= 8'b00000000;
		ins[114] <= 8'b00000000;
		ins[115] <= 8'b00000000;
	end

	assign ins_out = {ins[address + 3], ins[address + 2], ins[address + 1], ins[address]};
endmodule
